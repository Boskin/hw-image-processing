module vga640_480(

);

endmodule
